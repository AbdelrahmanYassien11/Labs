package simpleadder_pkg;

	`include "transaction.svh"

	`include "driver.svh"
	`include "inputMonitor.svh"
	`include "outputMonitor.svh"

	`include "predictor.svh"
	`include "comparator.svh"
	`include "scoreboard.svh"
	
	`include "randomized_sequence.svh"
	`include "test.svh"


endpackage